module a10_mac_8bitx2 (
		input  wire        clock0,  //  clock0.clock0
		input  wire [7:0]  dataa_0, // dataa_0.dataa_0
		input  wire [7:0]  dataa_1, // dataa_1.dataa_1
		input  wire [7:0]  datab_0, // datab_0.datab_0
		input  wire [7:0]  datab_1, // datab_1.datab_1
		output wire [31:0] result   //  result.result
	);
endmodule

